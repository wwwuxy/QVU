/* verilator lint_off WIDTHEXPAND */
module verilator_directives;
  // 空模块，仅用于添加Verilator属性
endmodule
/* verilator lint_on WIDTHEXPAND */
